
module niosv (
	clk_50m_clk,
	key_export,
	led_export,
	reset_50m_reset_n);	

	input		clk_50m_clk;
	input		key_export;
	output		led_export;
	input		reset_50m_reset_n;
endmodule
