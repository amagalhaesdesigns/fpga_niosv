-- niosv.vhd

-- Generated using ACDS version 23.1 991

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity niosv is
	port (
		clk_50m_clk       : in  std_logic := '0'; --   clk_50m.clk
		key_export        : in  std_logic := '0'; --       key.export
		led_export        : out std_logic;        --       led.export
		reset_50m_reset_n : in  std_logic := '0'  -- reset_50m.reset_n
	);
end entity niosv;

architecture rtl of niosv is
	component niosv_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component niosv_jtag_uart;

	component niosv_key is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component niosv_key;

	component niosv_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component niosv_led;

	component niosv_niosv is
		port (
			clk                          : in  std_logic                     := 'X';             -- clk
			reset_reset                  : in  std_logic                     := 'X';             -- reset
			platform_irq_rx_irq          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- irq
			instruction_manager_awaddr   : out std_logic_vector(31 downto 0);                    -- awaddr
			instruction_manager_awsize   : out std_logic_vector(2 downto 0);                     -- awsize
			instruction_manager_awlen    : out std_logic_vector(7 downto 0);                     -- awlen
			instruction_manager_awprot   : out std_logic_vector(2 downto 0);                     -- awprot
			instruction_manager_awvalid  : out std_logic;                                        -- awvalid
			instruction_manager_awburst  : out std_logic_vector(1 downto 0);                     -- awburst
			instruction_manager_awready  : in  std_logic                     := 'X';             -- awready
			instruction_manager_wdata    : out std_logic_vector(31 downto 0);                    -- wdata
			instruction_manager_wstrb    : out std_logic_vector(3 downto 0);                     -- wstrb
			instruction_manager_wlast    : out std_logic;                                        -- wlast
			instruction_manager_wvalid   : out std_logic;                                        -- wvalid
			instruction_manager_wready   : in  std_logic                     := 'X';             -- wready
			instruction_manager_bresp    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			instruction_manager_bvalid   : in  std_logic                     := 'X';             -- bvalid
			instruction_manager_bready   : out std_logic;                                        -- bready
			instruction_manager_araddr   : out std_logic_vector(31 downto 0);                    -- araddr
			instruction_manager_arsize   : out std_logic_vector(2 downto 0);                     -- arsize
			instruction_manager_arlen    : out std_logic_vector(7 downto 0);                     -- arlen
			instruction_manager_arprot   : out std_logic_vector(2 downto 0);                     -- arprot
			instruction_manager_arvalid  : out std_logic;                                        -- arvalid
			instruction_manager_arburst  : out std_logic_vector(1 downto 0);                     -- arburst
			instruction_manager_arready  : in  std_logic                     := 'X';             -- arready
			instruction_manager_rdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			instruction_manager_rresp    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			instruction_manager_rvalid   : in  std_logic                     := 'X';             -- rvalid
			instruction_manager_rready   : out std_logic;                                        -- rready
			instruction_manager_rlast    : in  std_logic                     := 'X';             -- rlast
			data_manager_awaddr          : out std_logic_vector(31 downto 0);                    -- awaddr
			data_manager_awsize          : out std_logic_vector(2 downto 0);                     -- awsize
			data_manager_awlen           : out std_logic_vector(7 downto 0);                     -- awlen
			data_manager_awprot          : out std_logic_vector(2 downto 0);                     -- awprot
			data_manager_awvalid         : out std_logic;                                        -- awvalid
			data_manager_awready         : in  std_logic                     := 'X';             -- awready
			data_manager_wdata           : out std_logic_vector(31 downto 0);                    -- wdata
			data_manager_wstrb           : out std_logic_vector(3 downto 0);                     -- wstrb
			data_manager_wlast           : out std_logic;                                        -- wlast
			data_manager_wvalid          : out std_logic;                                        -- wvalid
			data_manager_wready          : in  std_logic                     := 'X';             -- wready
			data_manager_bresp           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			data_manager_bvalid          : in  std_logic                     := 'X';             -- bvalid
			data_manager_bready          : out std_logic;                                        -- bready
			data_manager_araddr          : out std_logic_vector(31 downto 0);                    -- araddr
			data_manager_arsize          : out std_logic_vector(2 downto 0);                     -- arsize
			data_manager_arlen           : out std_logic_vector(7 downto 0);                     -- arlen
			data_manager_arprot          : out std_logic_vector(2 downto 0);                     -- arprot
			data_manager_arvalid         : out std_logic;                                        -- arvalid
			data_manager_arready         : in  std_logic                     := 'X';             -- arready
			data_manager_rdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			data_manager_rresp           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			data_manager_rvalid          : in  std_logic                     := 'X';             -- rvalid
			data_manager_rlast           : in  std_logic                     := 'X';             -- rlast
			data_manager_rready          : out std_logic;                                        -- rready
			ndm_reset_in_reset           : in  std_logic                     := 'X';             -- reset
			timer_sw_agent_write         : in  std_logic                     := 'X';             -- write
			timer_sw_agent_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			timer_sw_agent_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			timer_sw_agent_address       : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			timer_sw_agent_read          : in  std_logic                     := 'X';             -- read
			timer_sw_agent_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			timer_sw_agent_readdatavalid : out std_logic;                                        -- readdatavalid
			timer_sw_agent_waitrequest   : out std_logic;                                        -- waitrequest
			dm_agent_write               : in  std_logic                     := 'X';             -- write
			dm_agent_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dm_agent_address             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			dm_agent_read                : in  std_logic                     := 'X';             -- read
			dm_agent_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			dm_agent_readdatavalid       : out std_logic;                                        -- readdatavalid
			dm_agent_waitrequest         : out std_logic;                                        -- waitrequest
			dbg_reset_out_reset          : out std_logic                                         -- reset
		);
	end component niosv_niosv;

	component niosv_onchip_memory2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component niosv_onchip_memory2;

	component niosv_sys_clk is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component niosv_sys_clk;

	component niosv_mm_interconnect_0 is
		port (
			niosv_data_manager_awaddr                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			niosv_data_manager_awlen                    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- awlen
			niosv_data_manager_awsize                   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			niosv_data_manager_awprot                   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			niosv_data_manager_awvalid                  : in  std_logic                     := 'X';             -- awvalid
			niosv_data_manager_awready                  : out std_logic;                                        -- awready
			niosv_data_manager_wdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			niosv_data_manager_wstrb                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			niosv_data_manager_wlast                    : in  std_logic                     := 'X';             -- wlast
			niosv_data_manager_wvalid                   : in  std_logic                     := 'X';             -- wvalid
			niosv_data_manager_wready                   : out std_logic;                                        -- wready
			niosv_data_manager_bresp                    : out std_logic_vector(1 downto 0);                     -- bresp
			niosv_data_manager_bvalid                   : out std_logic;                                        -- bvalid
			niosv_data_manager_bready                   : in  std_logic                     := 'X';             -- bready
			niosv_data_manager_araddr                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			niosv_data_manager_arlen                    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- arlen
			niosv_data_manager_arsize                   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			niosv_data_manager_arprot                   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			niosv_data_manager_arvalid                  : in  std_logic                     := 'X';             -- arvalid
			niosv_data_manager_arready                  : out std_logic;                                        -- arready
			niosv_data_manager_rdata                    : out std_logic_vector(31 downto 0);                    -- rdata
			niosv_data_manager_rresp                    : out std_logic_vector(1 downto 0);                     -- rresp
			niosv_data_manager_rlast                    : out std_logic;                                        -- rlast
			niosv_data_manager_rvalid                   : out std_logic;                                        -- rvalid
			niosv_data_manager_rready                   : in  std_logic                     := 'X';             -- rready
			niosv_instruction_manager_awaddr            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			niosv_instruction_manager_awlen             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- awlen
			niosv_instruction_manager_awsize            : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			niosv_instruction_manager_awburst           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			niosv_instruction_manager_awprot            : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			niosv_instruction_manager_awvalid           : in  std_logic                     := 'X';             -- awvalid
			niosv_instruction_manager_awready           : out std_logic;                                        -- awready
			niosv_instruction_manager_wdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			niosv_instruction_manager_wstrb             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			niosv_instruction_manager_wlast             : in  std_logic                     := 'X';             -- wlast
			niosv_instruction_manager_wvalid            : in  std_logic                     := 'X';             -- wvalid
			niosv_instruction_manager_wready            : out std_logic;                                        -- wready
			niosv_instruction_manager_bresp             : out std_logic_vector(1 downto 0);                     -- bresp
			niosv_instruction_manager_bvalid            : out std_logic;                                        -- bvalid
			niosv_instruction_manager_bready            : in  std_logic                     := 'X';             -- bready
			niosv_instruction_manager_araddr            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			niosv_instruction_manager_arlen             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- arlen
			niosv_instruction_manager_arsize            : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			niosv_instruction_manager_arburst           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			niosv_instruction_manager_arprot            : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			niosv_instruction_manager_arvalid           : in  std_logic                     := 'X';             -- arvalid
			niosv_instruction_manager_arready           : out std_logic;                                        -- arready
			niosv_instruction_manager_rdata             : out std_logic_vector(31 downto 0);                    -- rdata
			niosv_instruction_manager_rresp             : out std_logic_vector(1 downto 0);                     -- rresp
			niosv_instruction_manager_rlast             : out std_logic;                                        -- rlast
			niosv_instruction_manager_rvalid            : out std_logic;                                        -- rvalid
			niosv_instruction_manager_rready            : in  std_logic                     := 'X';             -- rready
			clk_50m_clk_clk                             : in  std_logic                     := 'X';             -- clk
			jtag_uart_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			niosv_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			jtag_uart_avalon_jtag_slave_address         : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write           : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read            : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata       : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest     : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect      : out std_logic;                                        -- chipselect
			key_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			key_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_s1_address                              : out std_logic_vector(2 downto 0);                     -- address
			led_s1_write                                : out std_logic;                                        -- write
			led_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			led_s1_chipselect                           : out std_logic;                                        -- chipselect
			niosv_dm_agent_address                      : out std_logic_vector(15 downto 0);                    -- address
			niosv_dm_agent_write                        : out std_logic;                                        -- write
			niosv_dm_agent_read                         : out std_logic;                                        -- read
			niosv_dm_agent_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			niosv_dm_agent_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			niosv_dm_agent_readdatavalid                : in  std_logic                     := 'X';             -- readdatavalid
			niosv_dm_agent_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			niosv_timer_sw_agent_address                : out std_logic_vector(5 downto 0);                     -- address
			niosv_timer_sw_agent_write                  : out std_logic;                                        -- write
			niosv_timer_sw_agent_read                   : out std_logic;                                        -- read
			niosv_timer_sw_agent_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			niosv_timer_sw_agent_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			niosv_timer_sw_agent_byteenable             : out std_logic_vector(3 downto 0);                     -- byteenable
			niosv_timer_sw_agent_readdatavalid          : in  std_logic                     := 'X';             -- readdatavalid
			niosv_timer_sw_agent_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			onchip_memory2_s1_address                   : out std_logic_vector(15 downto 0);                    -- address
			onchip_memory2_s1_write                     : out std_logic;                                        -- write
			onchip_memory2_s1_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_s1_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_s1_byteenable                : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_s1_chipselect                : out std_logic;                                        -- chipselect
			onchip_memory2_s1_clken                     : out std_logic;                                        -- clken
			sys_clk_s1_address                          : out std_logic_vector(2 downto 0);                     -- address
			sys_clk_s1_write                            : out std_logic;                                        -- write
			sys_clk_s1_readdata                         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_clk_s1_writedata                        : out std_logic_vector(15 downto 0);                    -- writedata
			sys_clk_s1_chipselect                       : out std_logic                                         -- chipselect
		);
	end component niosv_mm_interconnect_0;

	component niosv_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(15 downto 0)         -- irq
		);
	end component niosv_irq_mapper;

	component niosv_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component niosv_rst_controller;

	component niosv_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component niosv_rst_controller_001;

	signal niosv_data_manager_arlen                                      : std_logic_vector(7 downto 0);  -- niosv:data_manager_arlen -> mm_interconnect_0:niosv_data_manager_arlen
	signal niosv_data_manager_wstrb                                      : std_logic_vector(3 downto 0);  -- niosv:data_manager_wstrb -> mm_interconnect_0:niosv_data_manager_wstrb
	signal niosv_data_manager_wready                                     : std_logic;                     -- mm_interconnect_0:niosv_data_manager_wready -> niosv:data_manager_wready
	signal niosv_data_manager_rready                                     : std_logic;                     -- niosv:data_manager_rready -> mm_interconnect_0:niosv_data_manager_rready
	signal niosv_data_manager_awlen                                      : std_logic_vector(7 downto 0);  -- niosv:data_manager_awlen -> mm_interconnect_0:niosv_data_manager_awlen
	signal niosv_data_manager_wvalid                                     : std_logic;                     -- niosv:data_manager_wvalid -> mm_interconnect_0:niosv_data_manager_wvalid
	signal niosv_data_manager_araddr                                     : std_logic_vector(31 downto 0); -- niosv:data_manager_araddr -> mm_interconnect_0:niosv_data_manager_araddr
	signal niosv_data_manager_arprot                                     : std_logic_vector(2 downto 0);  -- niosv:data_manager_arprot -> mm_interconnect_0:niosv_data_manager_arprot
	signal niosv_data_manager_awprot                                     : std_logic_vector(2 downto 0);  -- niosv:data_manager_awprot -> mm_interconnect_0:niosv_data_manager_awprot
	signal niosv_data_manager_wdata                                      : std_logic_vector(31 downto 0); -- niosv:data_manager_wdata -> mm_interconnect_0:niosv_data_manager_wdata
	signal niosv_data_manager_arvalid                                    : std_logic;                     -- niosv:data_manager_arvalid -> mm_interconnect_0:niosv_data_manager_arvalid
	signal niosv_data_manager_awaddr                                     : std_logic_vector(31 downto 0); -- niosv:data_manager_awaddr -> mm_interconnect_0:niosv_data_manager_awaddr
	signal niosv_data_manager_bresp                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:niosv_data_manager_bresp -> niosv:data_manager_bresp
	signal niosv_data_manager_arready                                    : std_logic;                     -- mm_interconnect_0:niosv_data_manager_arready -> niosv:data_manager_arready
	signal niosv_data_manager_rdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:niosv_data_manager_rdata -> niosv:data_manager_rdata
	signal niosv_data_manager_awready                                    : std_logic;                     -- mm_interconnect_0:niosv_data_manager_awready -> niosv:data_manager_awready
	signal niosv_data_manager_arsize                                     : std_logic_vector(2 downto 0);  -- niosv:data_manager_arsize -> mm_interconnect_0:niosv_data_manager_arsize
	signal niosv_data_manager_bready                                     : std_logic;                     -- niosv:data_manager_bready -> mm_interconnect_0:niosv_data_manager_bready
	signal niosv_data_manager_rlast                                      : std_logic;                     -- mm_interconnect_0:niosv_data_manager_rlast -> niosv:data_manager_rlast
	signal niosv_data_manager_wlast                                      : std_logic;                     -- niosv:data_manager_wlast -> mm_interconnect_0:niosv_data_manager_wlast
	signal niosv_data_manager_rresp                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:niosv_data_manager_rresp -> niosv:data_manager_rresp
	signal niosv_data_manager_bvalid                                     : std_logic;                     -- mm_interconnect_0:niosv_data_manager_bvalid -> niosv:data_manager_bvalid
	signal niosv_data_manager_awsize                                     : std_logic_vector(2 downto 0);  -- niosv:data_manager_awsize -> mm_interconnect_0:niosv_data_manager_awsize
	signal niosv_data_manager_awvalid                                    : std_logic;                     -- niosv:data_manager_awvalid -> mm_interconnect_0:niosv_data_manager_awvalid
	signal niosv_data_manager_rvalid                                     : std_logic;                     -- mm_interconnect_0:niosv_data_manager_rvalid -> niosv:data_manager_rvalid
	signal niosv_instruction_manager_awburst                             : std_logic_vector(1 downto 0);  -- niosv:instruction_manager_awburst -> mm_interconnect_0:niosv_instruction_manager_awburst
	signal niosv_instruction_manager_arlen                               : std_logic_vector(7 downto 0);  -- niosv:instruction_manager_arlen -> mm_interconnect_0:niosv_instruction_manager_arlen
	signal niosv_instruction_manager_wstrb                               : std_logic_vector(3 downto 0);  -- niosv:instruction_manager_wstrb -> mm_interconnect_0:niosv_instruction_manager_wstrb
	signal niosv_instruction_manager_wready                              : std_logic;                     -- mm_interconnect_0:niosv_instruction_manager_wready -> niosv:instruction_manager_wready
	signal niosv_instruction_manager_rready                              : std_logic;                     -- niosv:instruction_manager_rready -> mm_interconnect_0:niosv_instruction_manager_rready
	signal niosv_instruction_manager_awlen                               : std_logic_vector(7 downto 0);  -- niosv:instruction_manager_awlen -> mm_interconnect_0:niosv_instruction_manager_awlen
	signal niosv_instruction_manager_wvalid                              : std_logic;                     -- niosv:instruction_manager_wvalid -> mm_interconnect_0:niosv_instruction_manager_wvalid
	signal niosv_instruction_manager_araddr                              : std_logic_vector(31 downto 0); -- niosv:instruction_manager_araddr -> mm_interconnect_0:niosv_instruction_manager_araddr
	signal niosv_instruction_manager_arprot                              : std_logic_vector(2 downto 0);  -- niosv:instruction_manager_arprot -> mm_interconnect_0:niosv_instruction_manager_arprot
	signal niosv_instruction_manager_awprot                              : std_logic_vector(2 downto 0);  -- niosv:instruction_manager_awprot -> mm_interconnect_0:niosv_instruction_manager_awprot
	signal niosv_instruction_manager_wdata                               : std_logic_vector(31 downto 0); -- niosv:instruction_manager_wdata -> mm_interconnect_0:niosv_instruction_manager_wdata
	signal niosv_instruction_manager_arvalid                             : std_logic;                     -- niosv:instruction_manager_arvalid -> mm_interconnect_0:niosv_instruction_manager_arvalid
	signal niosv_instruction_manager_awaddr                              : std_logic_vector(31 downto 0); -- niosv:instruction_manager_awaddr -> mm_interconnect_0:niosv_instruction_manager_awaddr
	signal niosv_instruction_manager_bresp                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:niosv_instruction_manager_bresp -> niosv:instruction_manager_bresp
	signal niosv_instruction_manager_arready                             : std_logic;                     -- mm_interconnect_0:niosv_instruction_manager_arready -> niosv:instruction_manager_arready
	signal niosv_instruction_manager_rdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:niosv_instruction_manager_rdata -> niosv:instruction_manager_rdata
	signal niosv_instruction_manager_awready                             : std_logic;                     -- mm_interconnect_0:niosv_instruction_manager_awready -> niosv:instruction_manager_awready
	signal niosv_instruction_manager_arburst                             : std_logic_vector(1 downto 0);  -- niosv:instruction_manager_arburst -> mm_interconnect_0:niosv_instruction_manager_arburst
	signal niosv_instruction_manager_arsize                              : std_logic_vector(2 downto 0);  -- niosv:instruction_manager_arsize -> mm_interconnect_0:niosv_instruction_manager_arsize
	signal niosv_instruction_manager_bready                              : std_logic;                     -- niosv:instruction_manager_bready -> mm_interconnect_0:niosv_instruction_manager_bready
	signal niosv_instruction_manager_rlast                               : std_logic;                     -- mm_interconnect_0:niosv_instruction_manager_rlast -> niosv:instruction_manager_rlast
	signal niosv_instruction_manager_wlast                               : std_logic;                     -- niosv:instruction_manager_wlast -> mm_interconnect_0:niosv_instruction_manager_wlast
	signal niosv_instruction_manager_rresp                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:niosv_instruction_manager_rresp -> niosv:instruction_manager_rresp
	signal niosv_instruction_manager_bvalid                              : std_logic;                     -- mm_interconnect_0:niosv_instruction_manager_bvalid -> niosv:instruction_manager_bvalid
	signal niosv_instruction_manager_awsize                              : std_logic_vector(2 downto 0);  -- niosv:instruction_manager_awsize -> mm_interconnect_0:niosv_instruction_manager_awsize
	signal niosv_instruction_manager_awvalid                             : std_logic;                     -- niosv:instruction_manager_awvalid -> mm_interconnect_0:niosv_instruction_manager_awvalid
	signal niosv_instruction_manager_rvalid                              : std_logic;                     -- mm_interconnect_0:niosv_instruction_manager_rvalid -> niosv:instruction_manager_rvalid
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_niosv_dm_agent_readdata                     : std_logic_vector(31 downto 0); -- niosv:dm_agent_readdata -> mm_interconnect_0:niosv_dm_agent_readdata
	signal mm_interconnect_0_niosv_dm_agent_waitrequest                  : std_logic;                     -- niosv:dm_agent_waitrequest -> mm_interconnect_0:niosv_dm_agent_waitrequest
	signal mm_interconnect_0_niosv_dm_agent_address                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:niosv_dm_agent_address -> niosv:dm_agent_address
	signal mm_interconnect_0_niosv_dm_agent_read                         : std_logic;                     -- mm_interconnect_0:niosv_dm_agent_read -> niosv:dm_agent_read
	signal mm_interconnect_0_niosv_dm_agent_readdatavalid                : std_logic;                     -- niosv:dm_agent_readdatavalid -> mm_interconnect_0:niosv_dm_agent_readdatavalid
	signal mm_interconnect_0_niosv_dm_agent_write                        : std_logic;                     -- mm_interconnect_0:niosv_dm_agent_write -> niosv:dm_agent_write
	signal mm_interconnect_0_niosv_dm_agent_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:niosv_dm_agent_writedata -> niosv:dm_agent_writedata
	signal mm_interconnect_0_onchip_memory2_s1_chipselect                : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	signal mm_interconnect_0_onchip_memory2_s1_readdata                  : std_logic_vector(31 downto 0); -- onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	signal mm_interconnect_0_onchip_memory2_s1_address                   : std_logic_vector(15 downto 0); -- mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	signal mm_interconnect_0_onchip_memory2_s1_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	signal mm_interconnect_0_onchip_memory2_s1_write                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	signal mm_interconnect_0_onchip_memory2_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	signal mm_interconnect_0_onchip_memory2_s1_clken                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	signal mm_interconnect_0_led_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:led_s1_chipselect -> led:chipselect
	signal mm_interconnect_0_led_s1_readdata                             : std_logic_vector(31 downto 0); -- led:readdata -> mm_interconnect_0:led_s1_readdata
	signal mm_interconnect_0_led_s1_address                              : std_logic_vector(2 downto 0);  -- mm_interconnect_0:led_s1_address -> led:address
	signal mm_interconnect_0_led_s1_write                                : std_logic;                     -- mm_interconnect_0:led_s1_write -> mm_interconnect_0_led_s1_write:in
	signal mm_interconnect_0_led_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_s1_writedata -> led:writedata
	signal mm_interconnect_0_key_s1_readdata                             : std_logic_vector(31 downto 0); -- key:readdata -> mm_interconnect_0:key_s1_readdata
	signal mm_interconnect_0_key_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:key_s1_address -> key:address
	signal mm_interconnect_0_sys_clk_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:sys_clk_s1_chipselect -> sys_clk:chipselect
	signal mm_interconnect_0_sys_clk_s1_readdata                         : std_logic_vector(15 downto 0); -- sys_clk:readdata -> mm_interconnect_0:sys_clk_s1_readdata
	signal mm_interconnect_0_sys_clk_s1_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:sys_clk_s1_address -> sys_clk:address
	signal mm_interconnect_0_sys_clk_s1_write                            : std_logic;                     -- mm_interconnect_0:sys_clk_s1_write -> mm_interconnect_0_sys_clk_s1_write:in
	signal mm_interconnect_0_sys_clk_s1_writedata                        : std_logic_vector(15 downto 0); -- mm_interconnect_0:sys_clk_s1_writedata -> sys_clk:writedata
	signal mm_interconnect_0_niosv_timer_sw_agent_readdata               : std_logic_vector(31 downto 0); -- niosv:timer_sw_agent_readdata -> mm_interconnect_0:niosv_timer_sw_agent_readdata
	signal mm_interconnect_0_niosv_timer_sw_agent_waitrequest            : std_logic;                     -- niosv:timer_sw_agent_waitrequest -> mm_interconnect_0:niosv_timer_sw_agent_waitrequest
	signal mm_interconnect_0_niosv_timer_sw_agent_address                : std_logic_vector(5 downto 0);  -- mm_interconnect_0:niosv_timer_sw_agent_address -> niosv:timer_sw_agent_address
	signal mm_interconnect_0_niosv_timer_sw_agent_read                   : std_logic;                     -- mm_interconnect_0:niosv_timer_sw_agent_read -> niosv:timer_sw_agent_read
	signal mm_interconnect_0_niosv_timer_sw_agent_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:niosv_timer_sw_agent_byteenable -> niosv:timer_sw_agent_byteenable
	signal mm_interconnect_0_niosv_timer_sw_agent_readdatavalid          : std_logic;                     -- niosv:timer_sw_agent_readdatavalid -> mm_interconnect_0:niosv_timer_sw_agent_readdatavalid
	signal mm_interconnect_0_niosv_timer_sw_agent_write                  : std_logic;                     -- mm_interconnect_0:niosv_timer_sw_agent_write -> niosv:timer_sw_agent_write
	signal mm_interconnect_0_niosv_timer_sw_agent_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:niosv_timer_sw_agent_writedata -> niosv:timer_sw_agent_writedata
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- sys_clk:irq -> irq_mapper:receiver1_irq
	signal niosv_platform_irq_rx_irq                                     : std_logic_vector(15 downto 0); -- irq_mapper:sender_irq -> niosv:platform_irq_rx_irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, niosv:ndm_reset_in_reset, onchip_memory2:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:niosv_reset_reset_bridge_in_reset_reset, niosv:reset_reset]
	signal niosv_dbg_reset_out_reset                                     : std_logic;                     -- niosv:dbg_reset_out_reset -> rst_controller_001:reset_in1
	signal reset_50m_reset_n_ports_inv                                   : std_logic;                     -- reset_50m_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_led_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_led_s1_write:inv -> led:write_n
	signal mm_interconnect_0_sys_clk_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_sys_clk_s1_write:inv -> sys_clk:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [jtag_uart:rst_n, key:reset_n, led:reset_n, sys_clk:reset_n]

begin

	jtag_uart : component niosv_jtag_uart
		port map (
			clk            => clk_50m_clk,                                                   --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	key : component niosv_key
		port map (
			clk      => clk_50m_clk,                              --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_key_s1_address,         --                  s1.address
			readdata => mm_interconnect_0_key_s1_readdata,        --                    .readdata
			in_port  => key_export                                -- external_connection.export
		);

	led : component niosv_led
		port map (
			clk        => clk_50m_clk,                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_s1_readdata,        --                    .readdata
			out_port   => led_export                                -- external_connection.export
		);

	niosv : component niosv_niosv
		port map (
			clk                          => clk_50m_clk,                                          --                 clk.clk
			reset_reset                  => rst_controller_001_reset_out_reset,                   --               reset.reset
			platform_irq_rx_irq          => niosv_platform_irq_rx_irq,                            --     platform_irq_rx.irq
			instruction_manager_awaddr   => niosv_instruction_manager_awaddr,                     -- instruction_manager.awaddr
			instruction_manager_awsize   => niosv_instruction_manager_awsize,                     --                    .awsize
			instruction_manager_awlen    => niosv_instruction_manager_awlen,                      --                    .awlen
			instruction_manager_awprot   => niosv_instruction_manager_awprot,                     --                    .awprot
			instruction_manager_awvalid  => niosv_instruction_manager_awvalid,                    --                    .awvalid
			instruction_manager_awburst  => niosv_instruction_manager_awburst,                    --                    .awburst
			instruction_manager_awready  => niosv_instruction_manager_awready,                    --                    .awready
			instruction_manager_wdata    => niosv_instruction_manager_wdata,                      --                    .wdata
			instruction_manager_wstrb    => niosv_instruction_manager_wstrb,                      --                    .wstrb
			instruction_manager_wlast    => niosv_instruction_manager_wlast,                      --                    .wlast
			instruction_manager_wvalid   => niosv_instruction_manager_wvalid,                     --                    .wvalid
			instruction_manager_wready   => niosv_instruction_manager_wready,                     --                    .wready
			instruction_manager_bresp    => niosv_instruction_manager_bresp,                      --                    .bresp
			instruction_manager_bvalid   => niosv_instruction_manager_bvalid,                     --                    .bvalid
			instruction_manager_bready   => niosv_instruction_manager_bready,                     --                    .bready
			instruction_manager_araddr   => niosv_instruction_manager_araddr,                     --                    .araddr
			instruction_manager_arsize   => niosv_instruction_manager_arsize,                     --                    .arsize
			instruction_manager_arlen    => niosv_instruction_manager_arlen,                      --                    .arlen
			instruction_manager_arprot   => niosv_instruction_manager_arprot,                     --                    .arprot
			instruction_manager_arvalid  => niosv_instruction_manager_arvalid,                    --                    .arvalid
			instruction_manager_arburst  => niosv_instruction_manager_arburst,                    --                    .arburst
			instruction_manager_arready  => niosv_instruction_manager_arready,                    --                    .arready
			instruction_manager_rdata    => niosv_instruction_manager_rdata,                      --                    .rdata
			instruction_manager_rresp    => niosv_instruction_manager_rresp,                      --                    .rresp
			instruction_manager_rvalid   => niosv_instruction_manager_rvalid,                     --                    .rvalid
			instruction_manager_rready   => niosv_instruction_manager_rready,                     --                    .rready
			instruction_manager_rlast    => niosv_instruction_manager_rlast,                      --                    .rlast
			data_manager_awaddr          => niosv_data_manager_awaddr,                            --        data_manager.awaddr
			data_manager_awsize          => niosv_data_manager_awsize,                            --                    .awsize
			data_manager_awlen           => niosv_data_manager_awlen,                             --                    .awlen
			data_manager_awprot          => niosv_data_manager_awprot,                            --                    .awprot
			data_manager_awvalid         => niosv_data_manager_awvalid,                           --                    .awvalid
			data_manager_awready         => niosv_data_manager_awready,                           --                    .awready
			data_manager_wdata           => niosv_data_manager_wdata,                             --                    .wdata
			data_manager_wstrb           => niosv_data_manager_wstrb,                             --                    .wstrb
			data_manager_wlast           => niosv_data_manager_wlast,                             --                    .wlast
			data_manager_wvalid          => niosv_data_manager_wvalid,                            --                    .wvalid
			data_manager_wready          => niosv_data_manager_wready,                            --                    .wready
			data_manager_bresp           => niosv_data_manager_bresp,                             --                    .bresp
			data_manager_bvalid          => niosv_data_manager_bvalid,                            --                    .bvalid
			data_manager_bready          => niosv_data_manager_bready,                            --                    .bready
			data_manager_araddr          => niosv_data_manager_araddr,                            --                    .araddr
			data_manager_arsize          => niosv_data_manager_arsize,                            --                    .arsize
			data_manager_arlen           => niosv_data_manager_arlen,                             --                    .arlen
			data_manager_arprot          => niosv_data_manager_arprot,                            --                    .arprot
			data_manager_arvalid         => niosv_data_manager_arvalid,                           --                    .arvalid
			data_manager_arready         => niosv_data_manager_arready,                           --                    .arready
			data_manager_rdata           => niosv_data_manager_rdata,                             --                    .rdata
			data_manager_rresp           => niosv_data_manager_rresp,                             --                    .rresp
			data_manager_rvalid          => niosv_data_manager_rvalid,                            --                    .rvalid
			data_manager_rlast           => niosv_data_manager_rlast,                             --                    .rlast
			data_manager_rready          => niosv_data_manager_rready,                            --                    .rready
			ndm_reset_in_reset           => rst_controller_reset_out_reset,                       --        ndm_reset_in.reset
			timer_sw_agent_write         => mm_interconnect_0_niosv_timer_sw_agent_write,         --      timer_sw_agent.write
			timer_sw_agent_writedata     => mm_interconnect_0_niosv_timer_sw_agent_writedata,     --                    .writedata
			timer_sw_agent_byteenable    => mm_interconnect_0_niosv_timer_sw_agent_byteenable,    --                    .byteenable
			timer_sw_agent_address       => mm_interconnect_0_niosv_timer_sw_agent_address,       --                    .address
			timer_sw_agent_read          => mm_interconnect_0_niosv_timer_sw_agent_read,          --                    .read
			timer_sw_agent_readdata      => mm_interconnect_0_niosv_timer_sw_agent_readdata,      --                    .readdata
			timer_sw_agent_readdatavalid => mm_interconnect_0_niosv_timer_sw_agent_readdatavalid, --                    .readdatavalid
			timer_sw_agent_waitrequest   => mm_interconnect_0_niosv_timer_sw_agent_waitrequest,   --                    .waitrequest
			dm_agent_write               => mm_interconnect_0_niosv_dm_agent_write,               --            dm_agent.write
			dm_agent_writedata           => mm_interconnect_0_niosv_dm_agent_writedata,           --                    .writedata
			dm_agent_address             => mm_interconnect_0_niosv_dm_agent_address,             --                    .address
			dm_agent_read                => mm_interconnect_0_niosv_dm_agent_read,                --                    .read
			dm_agent_readdata            => mm_interconnect_0_niosv_dm_agent_readdata,            --                    .readdata
			dm_agent_readdatavalid       => mm_interconnect_0_niosv_dm_agent_readdatavalid,       --                    .readdatavalid
			dm_agent_waitrequest         => mm_interconnect_0_niosv_dm_agent_waitrequest,         --                    .waitrequest
			dbg_reset_out_reset          => niosv_dbg_reset_out_reset                             --       dbg_reset_out.reset
		);

	onchip_memory2 : component niosv_onchip_memory2
		port map (
			clk        => clk_50m_clk,                                    --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                 -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,             --       .reset_req
			freeze     => '0'                                             -- (terminated)
		);

	sys_clk : component niosv_sys_clk
		port map (
			clk        => clk_50m_clk,                                  --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_sys_clk_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_clk_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_clk_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_clk_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_clk_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                      --   irq.irq
		);

	mm_interconnect_0 : component niosv_mm_interconnect_0
		port map (
			niosv_data_manager_awaddr                   => niosv_data_manager_awaddr,                                 --                    niosv_data_manager.awaddr
			niosv_data_manager_awlen                    => niosv_data_manager_awlen,                                  --                                      .awlen
			niosv_data_manager_awsize                   => niosv_data_manager_awsize,                                 --                                      .awsize
			niosv_data_manager_awprot                   => niosv_data_manager_awprot,                                 --                                      .awprot
			niosv_data_manager_awvalid                  => niosv_data_manager_awvalid,                                --                                      .awvalid
			niosv_data_manager_awready                  => niosv_data_manager_awready,                                --                                      .awready
			niosv_data_manager_wdata                    => niosv_data_manager_wdata,                                  --                                      .wdata
			niosv_data_manager_wstrb                    => niosv_data_manager_wstrb,                                  --                                      .wstrb
			niosv_data_manager_wlast                    => niosv_data_manager_wlast,                                  --                                      .wlast
			niosv_data_manager_wvalid                   => niosv_data_manager_wvalid,                                 --                                      .wvalid
			niosv_data_manager_wready                   => niosv_data_manager_wready,                                 --                                      .wready
			niosv_data_manager_bresp                    => niosv_data_manager_bresp,                                  --                                      .bresp
			niosv_data_manager_bvalid                   => niosv_data_manager_bvalid,                                 --                                      .bvalid
			niosv_data_manager_bready                   => niosv_data_manager_bready,                                 --                                      .bready
			niosv_data_manager_araddr                   => niosv_data_manager_araddr,                                 --                                      .araddr
			niosv_data_manager_arlen                    => niosv_data_manager_arlen,                                  --                                      .arlen
			niosv_data_manager_arsize                   => niosv_data_manager_arsize,                                 --                                      .arsize
			niosv_data_manager_arprot                   => niosv_data_manager_arprot,                                 --                                      .arprot
			niosv_data_manager_arvalid                  => niosv_data_manager_arvalid,                                --                                      .arvalid
			niosv_data_manager_arready                  => niosv_data_manager_arready,                                --                                      .arready
			niosv_data_manager_rdata                    => niosv_data_manager_rdata,                                  --                                      .rdata
			niosv_data_manager_rresp                    => niosv_data_manager_rresp,                                  --                                      .rresp
			niosv_data_manager_rlast                    => niosv_data_manager_rlast,                                  --                                      .rlast
			niosv_data_manager_rvalid                   => niosv_data_manager_rvalid,                                 --                                      .rvalid
			niosv_data_manager_rready                   => niosv_data_manager_rready,                                 --                                      .rready
			niosv_instruction_manager_awaddr            => niosv_instruction_manager_awaddr,                          --             niosv_instruction_manager.awaddr
			niosv_instruction_manager_awlen             => niosv_instruction_manager_awlen,                           --                                      .awlen
			niosv_instruction_manager_awsize            => niosv_instruction_manager_awsize,                          --                                      .awsize
			niosv_instruction_manager_awburst           => niosv_instruction_manager_awburst,                         --                                      .awburst
			niosv_instruction_manager_awprot            => niosv_instruction_manager_awprot,                          --                                      .awprot
			niosv_instruction_manager_awvalid           => niosv_instruction_manager_awvalid,                         --                                      .awvalid
			niosv_instruction_manager_awready           => niosv_instruction_manager_awready,                         --                                      .awready
			niosv_instruction_manager_wdata             => niosv_instruction_manager_wdata,                           --                                      .wdata
			niosv_instruction_manager_wstrb             => niosv_instruction_manager_wstrb,                           --                                      .wstrb
			niosv_instruction_manager_wlast             => niosv_instruction_manager_wlast,                           --                                      .wlast
			niosv_instruction_manager_wvalid            => niosv_instruction_manager_wvalid,                          --                                      .wvalid
			niosv_instruction_manager_wready            => niosv_instruction_manager_wready,                          --                                      .wready
			niosv_instruction_manager_bresp             => niosv_instruction_manager_bresp,                           --                                      .bresp
			niosv_instruction_manager_bvalid            => niosv_instruction_manager_bvalid,                          --                                      .bvalid
			niosv_instruction_manager_bready            => niosv_instruction_manager_bready,                          --                                      .bready
			niosv_instruction_manager_araddr            => niosv_instruction_manager_araddr,                          --                                      .araddr
			niosv_instruction_manager_arlen             => niosv_instruction_manager_arlen,                           --                                      .arlen
			niosv_instruction_manager_arsize            => niosv_instruction_manager_arsize,                          --                                      .arsize
			niosv_instruction_manager_arburst           => niosv_instruction_manager_arburst,                         --                                      .arburst
			niosv_instruction_manager_arprot            => niosv_instruction_manager_arprot,                          --                                      .arprot
			niosv_instruction_manager_arvalid           => niosv_instruction_manager_arvalid,                         --                                      .arvalid
			niosv_instruction_manager_arready           => niosv_instruction_manager_arready,                         --                                      .arready
			niosv_instruction_manager_rdata             => niosv_instruction_manager_rdata,                           --                                      .rdata
			niosv_instruction_manager_rresp             => niosv_instruction_manager_rresp,                           --                                      .rresp
			niosv_instruction_manager_rlast             => niosv_instruction_manager_rlast,                           --                                      .rlast
			niosv_instruction_manager_rvalid            => niosv_instruction_manager_rvalid,                          --                                      .rvalid
			niosv_instruction_manager_rready            => niosv_instruction_manager_rready,                          --                                      .rready
			clk_50m_clk_clk                             => clk_50m_clk,                                               --                           clk_50m_clk.clk
			jtag_uart_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- jtag_uart_reset_reset_bridge_in_reset.reset
			niosv_reset_reset_bridge_in_reset_reset     => rst_controller_001_reset_out_reset,                        --     niosv_reset_reset_bridge_in_reset.reset
			jtag_uart_avalon_jtag_slave_address         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --           jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                      .write
			jtag_uart_avalon_jtag_slave_read            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                      .read
			jtag_uart_avalon_jtag_slave_readdata        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                      .readdata
			jtag_uart_avalon_jtag_slave_writedata       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                      .writedata
			jtag_uart_avalon_jtag_slave_waitrequest     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                      .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                      .chipselect
			key_s1_address                              => mm_interconnect_0_key_s1_address,                          --                                key_s1.address
			key_s1_readdata                             => mm_interconnect_0_key_s1_readdata,                         --                                      .readdata
			led_s1_address                              => mm_interconnect_0_led_s1_address,                          --                                led_s1.address
			led_s1_write                                => mm_interconnect_0_led_s1_write,                            --                                      .write
			led_s1_readdata                             => mm_interconnect_0_led_s1_readdata,                         --                                      .readdata
			led_s1_writedata                            => mm_interconnect_0_led_s1_writedata,                        --                                      .writedata
			led_s1_chipselect                           => mm_interconnect_0_led_s1_chipselect,                       --                                      .chipselect
			niosv_dm_agent_address                      => mm_interconnect_0_niosv_dm_agent_address,                  --                        niosv_dm_agent.address
			niosv_dm_agent_write                        => mm_interconnect_0_niosv_dm_agent_write,                    --                                      .write
			niosv_dm_agent_read                         => mm_interconnect_0_niosv_dm_agent_read,                     --                                      .read
			niosv_dm_agent_readdata                     => mm_interconnect_0_niosv_dm_agent_readdata,                 --                                      .readdata
			niosv_dm_agent_writedata                    => mm_interconnect_0_niosv_dm_agent_writedata,                --                                      .writedata
			niosv_dm_agent_readdatavalid                => mm_interconnect_0_niosv_dm_agent_readdatavalid,            --                                      .readdatavalid
			niosv_dm_agent_waitrequest                  => mm_interconnect_0_niosv_dm_agent_waitrequest,              --                                      .waitrequest
			niosv_timer_sw_agent_address                => mm_interconnect_0_niosv_timer_sw_agent_address,            --                  niosv_timer_sw_agent.address
			niosv_timer_sw_agent_write                  => mm_interconnect_0_niosv_timer_sw_agent_write,              --                                      .write
			niosv_timer_sw_agent_read                   => mm_interconnect_0_niosv_timer_sw_agent_read,               --                                      .read
			niosv_timer_sw_agent_readdata               => mm_interconnect_0_niosv_timer_sw_agent_readdata,           --                                      .readdata
			niosv_timer_sw_agent_writedata              => mm_interconnect_0_niosv_timer_sw_agent_writedata,          --                                      .writedata
			niosv_timer_sw_agent_byteenable             => mm_interconnect_0_niosv_timer_sw_agent_byteenable,         --                                      .byteenable
			niosv_timer_sw_agent_readdatavalid          => mm_interconnect_0_niosv_timer_sw_agent_readdatavalid,      --                                      .readdatavalid
			niosv_timer_sw_agent_waitrequest            => mm_interconnect_0_niosv_timer_sw_agent_waitrequest,        --                                      .waitrequest
			onchip_memory2_s1_address                   => mm_interconnect_0_onchip_memory2_s1_address,               --                     onchip_memory2_s1.address
			onchip_memory2_s1_write                     => mm_interconnect_0_onchip_memory2_s1_write,                 --                                      .write
			onchip_memory2_s1_readdata                  => mm_interconnect_0_onchip_memory2_s1_readdata,              --                                      .readdata
			onchip_memory2_s1_writedata                 => mm_interconnect_0_onchip_memory2_s1_writedata,             --                                      .writedata
			onchip_memory2_s1_byteenable                => mm_interconnect_0_onchip_memory2_s1_byteenable,            --                                      .byteenable
			onchip_memory2_s1_chipselect                => mm_interconnect_0_onchip_memory2_s1_chipselect,            --                                      .chipselect
			onchip_memory2_s1_clken                     => mm_interconnect_0_onchip_memory2_s1_clken,                 --                                      .clken
			sys_clk_s1_address                          => mm_interconnect_0_sys_clk_s1_address,                      --                            sys_clk_s1.address
			sys_clk_s1_write                            => mm_interconnect_0_sys_clk_s1_write,                        --                                      .write
			sys_clk_s1_readdata                         => mm_interconnect_0_sys_clk_s1_readdata,                     --                                      .readdata
			sys_clk_s1_writedata                        => mm_interconnect_0_sys_clk_s1_writedata,                    --                                      .writedata
			sys_clk_s1_chipselect                       => mm_interconnect_0_sys_clk_s1_chipselect                    --                                      .chipselect
		);

	irq_mapper : component niosv_irq_mapper
		port map (
			clk           => clk_50m_clk,                        --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			sender_irq    => niosv_platform_irq_rx_irq           --    sender.irq
		);

	rst_controller : component niosv_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_50m_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_50m_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component niosv_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_50m_reset_n_ports_inv,        -- reset_in0.reset
			reset_in1      => niosv_dbg_reset_out_reset,          -- reset_in1.reset
			clk            => clk_50m_clk,                        --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_50m_reset_n_ports_inv <= not reset_50m_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_led_s1_write_ports_inv <= not mm_interconnect_0_led_s1_write;

	mm_interconnect_0_sys_clk_s1_write_ports_inv <= not mm_interconnect_0_sys_clk_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of niosv
