-------------------------------------------------------------------------------
-- Title      : [Design Title, e.g., System Top Level]
-- Project    : [Project Name, e.g., Embedded Processor Projects]
-------------------------------------------------------------------------------
-- File       : fpga_niosv.vhd
-- Author     : Alexandre Magalhaes
-- Created    : September 29th, 2025
-- Last update: September 29th, 2025
-- Platform   : Intel/Altera Cyclone V]
-------------------------------------------------------------------------------
-- Description:
-- This template serves as the top-level entity for an FPGA design.
-- It is responsible for:
-- 1. Defining the primary I/O ports (clocks, resets, external interfaces).
-- 2. Instantiating and connecting internal system components (e.g., Nios V,
--    peripherals, custom logic).
--
-------------------------------------------------------------------------------

-- Libraries
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Top-level entity for the FPGA system.
entity fpga_niosv is
port (
    iClock      : in std_logic;  	-- The main input clock (e.g., 50 MHz).
    inReset     : in std_logic;  	-- The active-high or active-low system reset.
    iKey        : in std_logic;  	-- General purpose input (e.g., push-button).
    oLed        : out std_logic		-- General purpose output (e.g., status LED).
);
end entity;

architecture rtl of fpga_niosv is

    -- Internal signal declarations (e.g., clocks, resets, bus connections)
    -- signal internal_clock : std_logic;

    -- Component declaration for the Nios V processor.
    -- This component represents the design generated by Platform Designer (Qsys).
    component niosv is
        port (
            clk_50m_clk       : in  std_logic := 'X'; 	-- System Clock
            reset_50m_reset_n : in  std_logic := 'X';	-- Active-low Reset
            key_export        : in  std_logic := 'X'; 	-- Key input to the Nios V system
            led_export        : out std_logic        	-- LED output from the Nios V system
        );
    end component niosv;

begin

    -- Instance of the Nios V processor component.
    -- Map the top-level ports to the internal component ports.
    fpga_niosv_inst : component niosv
        port map (
            clk_50m_clk       => iClock,
            reset_50m_reset_n => inReset,
            key_export        => iKey,
            led_export        => oLed
        );
        
    -- Additional concurrent statements or processes for custom logic can be added here.
    
end architecture;